//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module parallel_to_serial
# (
    parameter width = 8
)
(
    input                      clk,
    input                      rst,

    input                      parallel_valid,
    input        [width - 1:0] parallel_data,

    output                     busy,
    output logic               serial_valid,
    output logic               serial_data
);
    // Task:
    // Implement a module that converts multi-bit parallel value to the single-bit serial data.
    //
    // The module should accept 'width' bit input parallel data when 'parallel_valid' input is asserted.
    // At the same clock cycle as 'parallel_valid' is asserted, the module should output
    // the least significant bit of the input data. In the following clock cycles the module
    // should output all the remaining bits of the parallel_data.
    // Together with providing correct 'serial_data' value, module should also assert the 'serial_valid' output.
    //
    // Note:
    // Check the waveform diagram in the README for better understanding.

    localparam w_index = $clog2 (width); 

    logic [w_index - 1:0] index = '0;
    logic [width - 1:0]reg_parallel_in_serial;

    always_ff @( posedge clk )
        
        if (rst)
            index <= '0;
        else
        begin
            if (parallel_valid)
                index <= 1'd1;
            else
            begin
                if (index > 1'd0) 
                begin

                    index <= index + 1'd1;
                    
                end
                else
                begin
                    
                    index <= '0;

                end
            end
        end
            

    always_ff @( posedge clk )     

        if (rst) 
        begin
            reg_parallel_in_serial <= '0;
        end 
        else 
        begin
            if (parallel_valid) 
            begin

                reg_parallel_in_serial <= parallel_data;

                
            end
        end

    //---------------------------------------------------- END BLOCK ----------------------------------------------------



    //---------------------------------------------------- OUTPUT SIGNALS -----------------------------------------------

    assign serial_valid  =  parallel_valid | index != w_index '(0);
    assign  serial_data  =  parallel_valid ? parallel_data[0] : reg_parallel_in_serial [index];
    assign         busy  =  index != w_index '(0) ? '1 : '0;




endmodule
