//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module sort_two_floats_ab (
    input        [FLEN - 1:0] a,
    input        [FLEN - 1:0] b,

    output logic [FLEN - 1:0] res0,
    output logic [FLEN - 1:0] res1,
    output                    err
);

    logic a_less_or_equal_b;

    f_less_or_equal i_floe (
        .a   ( a                 ),
        .b   ( b                 ),
        .res ( a_less_or_equal_b ),
        .err ( err               )
    );

    always_comb begin : a_b_compare
        if ( a_less_or_equal_b ) begin
            res0 = a;
            res1 = b;
        end
        else
        begin
            res0 = b;
            res1 = a;
        end
    end

endmodule

//----------------------------------------------------------------------------
// Example - different style
//----------------------------------------------------------------------------

module sort_two_floats_array
(
    input        [0:1][FLEN - 1:0] unsorted,
    output logic [0:1][FLEN - 1:0] sorted,
    output                         err
);

    logic u0_less_or_equal_u1;

    f_less_or_equal i_floe
    (
        .a   ( unsorted [0]        ),
        .b   ( unsorted [1]        ),
        .res ( u0_less_or_equal_u1 ),
        .err ( err                 )
    );

    always_comb
        if (u0_less_or_equal_u1)
            sorted = unsorted;
        else
              {   sorted [0],   sorted [1] }
            = { unsorted [1], unsorted [0] };

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module sort_three_floats (
    input        [0:2][FLEN - 1:0] unsorted,
    output logic [0:2][FLEN - 1:0] sorted,
    output                         err
);

    // Task:
    // Implement a module that accepts three Floating-Point numbers and outputs them in the increasing order.
    // The module should be combinational with zero latency.
    // The solution can use up to three instances of the "f_less_or_equal" module.
    //
    // Notes:
    // res0 must be less or equal to the res1
    // res1 must be less or equal to the res2
    //
    // The FLEN parameter is defined in the "import/preprocessed/cvw/config-shared.vh" file
    // and usually equal to the bit width of the double-precision floating-point number, FP64, 64 bits.

    logic u0_less_or_equal_u1, u1_less_or_equal_u2, u0_less_or_equal_u2;
    logic err_0_1, err_0_2, err_1_2;

    f_less_or_equal i_floe_0_1
    (
        .a   ( unsorted [0]        ), //a
        .b   ( unsorted [1]        ), //b
        .res ( u0_less_or_equal_u1 ),
        .err ( err_0_1             )
    );

    f_less_or_equal i_floe_1_2
    (
        .a   ( unsorted [1]        ), //b
        .b   ( unsorted [2]        ), //c
        .res ( u1_less_or_equal_u2 ),
        .err ( err_1_2             )
    );

    f_less_or_equal i_floe_0_2
    (
        .a   ( unsorted [0]        ), //a
        .b   ( unsorted [2]        ), //c
        .res ( u0_less_or_equal_u2 ),
        .err ( err_0_2             )
    );

    // a<b b<c, a<b<c
    // a<b b>c, a?c -> 1) a<c<b 2) c<a<b
    // a>b b<c, a?c -> 1) b<a<c 2) b<c<a
    // a>b b>c, c<b<a


    logic [0:2][FLEN - 1:0] mux_out;
    always_comb
    begin

        case ({u0_less_or_equal_u2,u1_less_or_equal_u2,u0_less_or_equal_u1}) // {a?c, b?c, a?b}
            3'b?11     :                            mux_out      =  unsorted                                  ; // a<b<c
            3'b101     : {mux_out [0], mux_out [1], mux_out [2]} = {unsorted [0], unsorted [2], unsorted [1]} ; // a<c<b
            3'b001     : {mux_out [0], mux_out [1], mux_out [2]} = {unsorted [2], unsorted [0], unsorted [1]} ; // c<a<b
            3'b110     : {mux_out [0], mux_out [1], mux_out [2]} = {unsorted [1], unsorted [0], unsorted [2]} ; // b<a<c
            3'b010     : {mux_out [0], mux_out [1], mux_out [2]} = {unsorted [1], unsorted [2], unsorted [0]} ; // b<c<a
            3'b000     : {mux_out [0], mux_out [1], mux_out [2]} = {unsorted [2], unsorted [1], unsorted [0]} ; // c<b<a
            default    :                            mux_out      =  unsorted                                  ;
        endcase
    end


    assign sorted = mux_out;
    assign err = |{err_0_2, err_1_2, err_0_1}; // Хотя бы один err

endmodule
